//conv build in 3*3*3 convlution core
//for 6*6*3 input data 

module CONV3 (
    input clk,
    input rst,
    input conv_en,
    output conv_done,
    input [7:0] conv_in,
    output [7:0] conv_out
);
    
endmodule