module moduleName (
  ports
);

endmodule
